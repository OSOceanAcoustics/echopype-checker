netcdf echopype-test-D20211005-T001612 {

// global attributes:
    :conventions = "CF-1.7, SONAR-netCDF4-1.0, ACDD-1.3" ;
    :keywords = "EK80" ;
    :sonar_convention_authority = "ICES" ;
    :sonar_convention_name = "SONAR-netCDF4" ;
    :sonar_convention_version = "1.0" ;
    :summary = "" ;
    :title = "" ;
    :date_created = "2021-10-05T00:16:12Z" ;
    :survey_name = "" ;

group: Environment {
  dimensions:
    time1 = 1 ;
    sound_velocity_profile_depth = 2 ;
   // missing frequency dimension
  variables:
    // missing frequency (M), absorption_indicative (M)
   // add long_name, standard_name and units to several variables
    double time1(time1) ;
      time1:_FillValue = NaN ;
      time1:axis = "T" ;
      time1:long_name = "Timestamps for NMEA position datagrams" ;
      time1:standard_name = "time" ;
      time1:comment = "Time coordinate corresponding to environmental variables. Note that Platform.time3 is the same as Environment.time1." ;
      time1:units = "seconds since 1900-01-01T00:00:00+00:00" ;
      time1:calendar = "gregorian" ;
      time1:echopype_mods = "added-allowed" ;
    double sound_velocity_profile_depth(sound_velocity_profile_depth) ;
      sound_velocity_profile_depth:_FillValue = NaN ;
      sound_velocity_profile_depth:standard_name = "depth" ;
      sound_velocity_profile_depth:units = "m" ;
      sound_velocity_profile_depth:axis = "Z" ;
      sound_velocity_profile_depth:positive = "down" ;
      sound_velocity_profile_depth:valid_min = 0. ;
      sound_velocity_profile_depth:echopype_mods = "added-allowed" ;
    float sound_speed_indicative(time1) ;
      sound_speed_indicative:long_name = "Indicative sound speed" ;
      sound_speed_indicative:standard_name = "speed_of_sound_in_sea_water" ;
      sound_speed_indicative:units = "m/s" ;
      sound_speed_indicative:valid_min = 0.0 ;
      sound_speed_indicative:_FillValue = NaN ;
   double depth(time1) ;
      depth:_FillValue = NaN ;
      depth:echopype_mods = "added-allowed" ;
    string transducer_name(time1) ;
      transducer_name:echopype_mods = "added-allowed" ;
    double transducer_sound_speed(time1) ;
      transducer_sound_speed:_FillValue = NaN ;
      transducer_sound_speed:echopype_mods = "added-allowed" ;
    double acidity(time1) ;
      acidity:_FillValue = NaN ;
      acidity:echopype_mods = "added-allowed" ;
    double salinity(time1) ;
      salinity:_FillValue = NaN ;
      salinity:echopype_mods = "added-allowed" ;
    double temperature(time1) ;
      temperature:_FillValue = NaN ;
      temperature:echopype_mods = "added-allowed" ;
    string sound_velocity_source(time1) ;
      sound_velocity_source:echopype_mods = "added-allowed" ;
    double sound_velocity_profile(time1, sound_velocity_profile_depth) ;
      sound_velocity_profile:long_name = "sound velocity profile" ;
      sound_velocity_profile:standard_name = "speed_of_sound_in_sea_water" ;
      sound_velocity_profile:units = "m/s" ;
      sound_velocity_profile:valid_min = 0. ;
      sound_velocity_profile:_FillValue = NaN ;
      sound_velocity_profile:comment = "parsed from raw data files as (depth, sound_speed) value pairs" ;
      sound_velocity_profile:echopype_mods = "added-allowed" ;
  data:

   depth = 100 ;

   acidity = 8 ;

   salinity = 35 ;

   temperature = 10 ;

   sound_speed_indicative = 1500 ;

   sound_velocity_profile = 1500, 1500 ;

   sound_velocity_source = "Calculated" ;

   transducer_name = "Unknown" ;

   transducer_sound_speed = 1500 ;

   time1 = 3842381772.962 ;

   sound_velocity_profile_depth = 1, 1000 ;
  } // group Environment

group: Platform {
  dimensions:
    channel = 3 ;
    time2 = 5 ;
    time1 = 1 ;
    time3 = 1 ;
  variables:
    // Not present: distance (O), heading (MA), speed_ground (MA), speed_relativ (O)
    double latitude(time1) ;
      latitude:_FillValue = NaN ;
      latitude:long_name = "Platform latitude" ;
      latitude:standard_name = "latitude" ;
      latitude:units = "degrees_north" ;
      latitude:valid_range = "(-90.0, 90.0)" ;
    double longitude(time1) ;
      longitude:_FillValue = NaN ;
      longitude:long_name = "Platform longitude" ;
      longitude:standard_name = "longitude" ;
      longitude:units = "degrees_east" ;
      longitude:valid_range = "(-180.0, 180.0)" ;
    uint64 time1(time1) ;
      time1:_FillValue = NaN ;
      time1:axis = "T" ;
      time1:long_name = "Timestamps for NMEA datagrams" ;
      time1:standard_name = "time" ;
      time1:comment = "Time coordinate corresponding to NMEA position data." ;
      time1:units = "seconds since 1900-01-01T00:00:00+00:00" ;
      time1:calendar = "gregorian" ;
    uint64 time2(time2) ;
      time2:_FillValue = NaN ;
      time2:axis = "T" ;
      time2:long_name = "Timestamps for platform motion and orientation data" ;
      time2:standard_name = "time" ;
      time2:comment = "Time coordinate corresponding to platform motion and orientation data." ;
      time2:units = "seconds since 1900-01-01T00:00:00+00:00" ;
      time2:calendar = "gregorian" ;
    uint64 time3(time3) ;
      time3:_FillValue = NaN ;
      time3:axis = "T" ;
      time3:long_name = "Timestamps for platform-related sampling environment" ;
      time3:standard_name = "time" ;
      time3:comment = "Time coordinate corresponding to platform-related sampling environment. Note that Platform.time3 is the same as Environment.time1." ;
      time3:units = "seconds since 1900-01-01T00:00:00+00:00" ;
      time3:calendar = "gregorian" ;
    string channel(channel) ;
      channel:long_name = "Vendor channel ID" ;
      channel:echopype_mods = "added" ;
   double frequency_nominal(channel) ;
      frequency_nominal:_FillValue = NaN ;
      frequency_nominal:units = "Hz" ;
      frequency_nominal:long_name = "Transducer frequency" ;
      frequency_nominal:valid_min = 0. ;
      frequency_nominal:standard_name = "sound_frequency" ;
      frequency_nominal:echopype_mods = "added" ;
    double pitch(time2) ;
      pitch:_FillValue = NaN ;
      pitch:long_name = "Platform pitch" ;
      pitch:standard_name = "platform_pitch_angle" ;
      pitch:units = "arc_degree" ;
      pitch:valid_range = "(-90.0, 90.0)" ;
    float roll(time2) ;
      roll:_FillValue = NaN ;
      roll:long_name = "Platform roll" ;
      roll:standard_name = "platform_roll_angle" ;
      roll:units = "arc_degree" ;
      roll:valid_range = "(-90.0, 90.0)" ; // valid range is supposed to be (-180.0, 180.0)
    float vertical_offset(time2) ;
      vertical_offset:_FillValue = NaN ;
      vertical_offset:long_name = "Platform vertical offset from nominal" ;
      vertical_offset:units = "m" ;
    float water_level(time3) ;
      water_level:_FillValue = NaN ;
      water_level:long_name = "z-axis distance from the platform coordinate system origin to the sonar transducer" ;
      water_level:units = "m" ;
    int64 water_level_draft_is_manual(time3) ;
      water_level_draft_is_manual:echopype_mods = "added" ;
    double sentence_type(time1) ;
      sentence_type:_FillValue = NaN ;
      sentence_type:echopype_mods = "added" ;
    double drop_keel_offset(time3) ;
      drop_keel_offset:_FillValue = NaN ;
      drop_keel_offset:echopype_mods = "added" ;
    int64 drop_keel_offset_is_manual(time3) ;
      drop_keel_offset_is_manual:echopype_mods = "added" ;
    float MRU_offset_x ;
      MRU_offset_x:_FillValue = NaN ;
      MRU_offset_x:long_name = "Distance along the x-axis from the platform coordinate system origin to the motion reference unit sensor origin" ;
      MRU_offset_x:units = "m" ;
    float MRU_offset_y ;
      MRU_offset_y:_FillValue = NaN ;
      MRU_offset_y:long_name = "Distance along the y-axis from the platform coordinate system origin to the motion reference unit sensor origin" ;
      MRU_offset_y:units = "m" ;
    float MRU_offset_z ;
      MRU_offset_z:_FillValue = NaN ;
      MRU_offset_z:long_name = "Distance along the z-axis from the platform coordinate system origin to the motion reference unit sensor origin" ;
      MRU_offset_z:units = "m" ;
    float MRU_rotation_x ;
      MRU_rotation_x:_FillValue = NaN ;
      MRU_rotation_x:long_name = "Extrinsic rotation about the x-axis from the platform to MRU coordinate systems" ;
      MRU_rotation_x:units = "arc_degree" ;
      MRU_rotation_x:valid_range = "(-180.0, 180.0)" ;
    float MRU_rotation_y ;
      MRU_rotation_y:_FillValue = NaN ;
      MRU_rotation_y:long_name = "Extrinsic rotation about the y-axis from the platform to MRU coordinate systems" ;
      MRU_rotation_y:units = "arc_degree" ;
      MRU_rotation_y:valid_range = "(-180.0, 180.0)" ;
    float MRU_rotation_z ;
      MRU_rotation_z:_FillValue = NaN ;
      MRU_rotation_z:long_name = "Extrinsic rotation about the z-axis from the platform to MRU coordinate systems" ;
      MRU_rotation_z:units = "arc_degree" ;
      MRU_rotation_z:valid_range = "(-180.0, 180.0)" ;
    float position_offset_x ;
      position_offset_x:_FillValue = NaN ;
      position_offset_x:long_name = "Distance along the x-axis from the platform coordinate system origin to the latitude/longitude sensor origin" ;
      position_offset_x:units = "m" ;
    float position_offset_y ;
      position_offset_y:_FillValue = NaN ;
      position_offset_y:long_name = "Distance along the y-axis from the platform coordinate system origin to the latitude/longitude sensor origin" ;
      position_offset_y:units = "m" ;
    float position_offset_z ;
      position_offset_z:_FillValue = NaN ;
      position_offset_z:long_name = "Distance along the z-axis from the platform coordinate system origin to the latitude/longitude sensor origin" ;
      position_offset_z:units = "m" ;
    float transducer_offset_x(channel) ;
      transducer_offset_x:_FillValue = NaN ;
      transducer_offset_x:long_name = "x-axis distance from the platform coordinate system origin to the sonar transducer" ;
      transducer_offset_x:units = "m" ;
    float transducer_offset_y(channel) ;
      transducer_offset_y:_FillValue = NaN ;
      transducer_offset_y:long_name = "y-axis distance from the platform coordinate system origin to the sonar transducer" ;
      transducer_offset_y:units = "m" ;
    float transducer_offset_z(channel) ;
      transducer_offset_z:_FillValue = NaN ;
      transducer_offset_z:long_name = "z-axis distance from the platform coordinate system origin to the sonar transducer" ;
      transducer_offset_z:units = "m" ;

  // group attributes:
      :platform_code_ICES = "" ;
      :platform_name = "" ;
      :platform_type = "" ;
  data:

   frequency_nominal = 120000, 200000, 70000 ;

   pitch = 0, 0, 0, 0, 0 ;

   roll = 0, 0, 0, 0, 0 ;

   vertical_offset = 0, 0, 0, 0, 0 ;

   latitude = _ ;

   longitude = _ ;

   sentence_type = _ ;

   drop_keel_offset = _ ;

   drop_keel_offset_is_manual = 0 ;

   transducer_offset_x = 0, 0, 0 ;

   transducer_offset_y = 0, 0, 0 ;

   transducer_offset_z = 0, 0, 0 ;

   water_level = 0 ;

   water_level_draft_is_manual = 0 ;

   MRU_offset_x = _ ;

   MRU_offset_y = _ ;

   MRU_offset_z = _ ;

   MRU_rotation_x = _ ;

   MRU_rotation_y = _ ;

   MRU_rotation_z = _ ;

   position_offset_x = _ ;

   position_offset_y = _ ;

   position_offset_z = _ ;

   channel = "WBT 150013-15 ES120-7C_ES", "WBT 545612-15 ES200-7C_ES", 
      "WBT 549762-15 ES70-7C_ES" ;

   time1 = _ ;

   time2 = 3842381772, 3842381773, 3842381774, 3842381775, 
      3842381776.964 ;

   time3 = 3842381772 ;


  group: NMEA {
    dimensions:
      // called "time" in convention
      time1 = 1 ;
    variables:
      string NMEA_datagram(time1) ;
        NMEA_datagram:long_name = "NMEA datagram" ;
      uint64 time1(time1) ;
        time1:_FillValue = NaN ;
        time1:axis = "T" ;
        time1:long_name = "Timestamps for NMEA datagrams" ;
        time1:standard_name = "time" ;
        time1:comment = "Time coordinate corresponding to NMEA sensor data." ;
        time1:units = "seconds since 1900-01-01T00:00:00+00:00" ;
        time1:calendar = "gregorian" ;
         time1:echopype_mods = "changed-attrs,changed-var" ;

    // group attributes:
        :description = "All NMEA sensor datagrams" ;
    data:

     NMEA_datagram = "$SDVLW,51.576,N,51.576,N" ;

     time1 = 3842381772 ;
    } // group NMEA
  } // group Platform

group: Provenance {
  dimensions:
    filenames = 1 ;
  variables:
    string source_filenames(filenames) ;
      source_filenames:long_name = "Source filenames" ;
    int64 filenames(filenames) ;
      filenames:long_name = "Index for data and metadata source filenames" ;

  // group attributes:
      :conversion_software_name = "echopype" ;
      :conversion_software_version = "0.6.4.dev112+g196bd6b2.d20230417" ;
      :conversion_time = "2023-05-18T03:39:38Z" ;
  data:

   source_filenames = "echopype-test-D20211005-T001612.raw" ;

   filenames = 0 ;
  } // group Provenance

group: Sonar {
  dimensions:
    channel = 3 ;
    beam_group = 2 ;
  variables:
    double frequency_nominal(channel) ;
      frequency_nominal:_FillValue = NaN ;
      frequency_nominal:units = "Hz" ;
      frequency_nominal:long_name = "Transducer frequency" ;
      frequency_nominal:valid_min = 0. ;
      frequency_nominal:standard_name = "sound_frequency" ;
      frequency_nominal:echopype_mods = "added" ;
    string channel(channel) ;
      channel:long_name = "Vendor channel ID" ;
      channel:echopype_mods = "added" ;
    string transceiver_serial_number(channel) ;
      transceiver_serial_number:long_name = "Transceiver serial number" ;
      transceiver_serial_number:echopype_mods = "added" ;
    string transducer_name(channel) ;
      transducer_name:long_name = "Transducer name" ;
      transducer_name:echopype_mods = "added" ;
    string transducer_serial_number(channel) ;
      transducer_serial_number:long_name = "Transducer serial number" ;
      :echopype_mods = "added" ;
    string beam_group(beam_group) ;
      beam_group:long_name = "Beam group name" ;
      beam_group:echopype_mods = "added" ;
    string beam_group_descr(beam_group) ;
      beam_group_descr:long_name = "Beam group description" ;
      beam_group_descr:echopype_mods = "added" ;

  // group attributes:
      :sonar_manufacturer = "Simrad" ;
      :sonar_model = "EK80" ;
      :sonar_serial_number = "" ;
      :sonar_software_name = "EK80" ;
      :sonar_software_version = "2.0.1.0" ;
      :sonar_type = "echosounder" ;
  data:

   frequency_nominal = 120000, 200000, 70000 ;

   transceiver_serial_number = "150013", "545612", "549762" ;

   transducer_name = "ES120-7C", "ES200-7C", "ES70-7C" ;

   transducer_serial_number = "1808", "213", "116" ;

   beam_group_descr = 
      "contains complex backscatter data and other beam or channel-specific data.", 
      "contains backscatter power (uncalibrated) and other beam or channel-specific data, including split-beam angle data when they exist." ;

   channel = "WBT 150013-15 ES120-7C_ES", "WBT 545612-15 ES200-7C_ES", 
      "WBT 549762-15 ES70-7C_ES" ;

   beam_group = "Beam_group1", "Beam_group2" ;

  group: Beam_group1 {
    dimensions:
      channel = 1 ;
      ping_time = 5 ;
      beam = 4 ;
      range_sample = 2 ;
    variables:
      // CONVENTION VARIABLES MISSING FROM EK80 IN ECHOPYPE
      // --- I have not modified the dimensions yet, nor added sample data or replaced use of enum types
      // Note: I've ommitted the beam_receive/transmit_minor/major variables.
      // Also ommitted MA variables described as necessary for type 1 and 2, 
      // (except for gain_correction and transmit_power):
      // receiver_sensitivity, time_varied_gain, transducer_gain, transmit_duration_equivalent, transmit_source_level
      beam_stabilisation_t beam_stabilisation(ping_time) ;
        beam_stabilisation:long_name =  "Beam stabilisation applied (or not)" ;
        beam_stabilisation:obligation = "M" ;
      float gain_correction(ping_time, beam) ;
        // This variable is found in EK60 and AZFP
        gain_correction:long_name = "Gain correction" ;
        gain_correction:units = "dB" ;
        gain_correction:obligation = "MA" ;
      short non_quantitative_processing(ping_time) ;
        non_quantitative_processing:flag_meanings = "strings" ;
        non_quantitative_processing:flag_values = 1,2 ;
        non_quantitative_processing:long_name = "Presence or not of non-quantitative processing applied to the backscattering data (sonar specific)" ;
        non_quantitative_processing:obligation = "M" ;
      float sample_time_offset(ping_time) ;
        sample_time_offset:long_name = "Time offset that is subtracted from the timestamp of each sample" ;
        sample_time_offset:units = "s" ;
        sample_time_offset:obligation = "M" ;
      float transmit_bandwidth(ping_time) ;
        transmit_bandwidth:long_name = "Nominal bandwidth of transmitted pulse" ;
        transmit_bandwidth:units = "Hz" ;
        transmit_bandwidth:valid_min = 0.0 ;
        transmit_bandwidth:obligation = "O" ;
      float transmit_frequency_start(ping_time, beam) ;
        transmit_frequency_start:long_name = "Start frequency in transmitted pulse" ;
        transmit_frequency_start:standard_name = "sound_frequency" ;
        transmit_frequency_start:units = "Hz" ;
        transmit_frequency_start:valid_min = 0.0 ;
        transmit_frequency_start:obligation = "M" ;
      float transmit_frequency_stop(ping_time, beam) ;
        transmit_frequency_stop:long_name = "Stop frequency in transmitted pulse" ;
        transmit_frequency_stop:standard_name = "sound_frequency" ;
        transmit_frequency_stop:units = "Hz" ;
        transmit_frequency_stop:valid_min = 0.0 ;
        transmit_frequency_stop:obligation = "M" ;
      transmit_t transmit_type(ping_time) ;
        transmit_type:long_name = "Type of transmitted pulse" ;
        transmit_type:obligation = "M" ;
      // ------------------------
      // ADDED FROM Beam_group2
      // Do they duplicate existing variables in Beam_group1?
      double angle_athwartship(channel, ping_time, range_sample, beam) ;
        angle_athwartship:_FillValue = NaN ;
        angle_athwartship:long_name = "electrical athwartship angle" ;
        angle_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
        :obligation = "NA" ;
        angle_athwartship:echopype_mods = "added" ;
      double angle_alongship(channel, ping_time, range_sample, beam) ;
        angle_alongship:_FillValue = NaN ;
        angle_alongship:long_name = "electrical alongship angle" ;
        angle_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
        :obligation = "NA" ;
        angle_alongship:echopype_mods = "added" ;
      // ------------------------
      double angle_offset_alongship(channel, ping_time, beam) ;
        angle_offset_alongship:_FillValue = NaN ;
        angle_offset_alongship:long_name = "electrical alongship angle offset of the transducer" ;
        angle_offset_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
        angle_offset_alongship:obligation = "NA" ;
        angle_offset_alongship:echopype_mods = "added" ;
      double angle_offset_athwartship(channel, ping_time, beam) ;
        angle_offset_athwartship:_FillValue = NaN ;
        angle_offset_athwartship:long_name = "electrical athwartship angle offset of the transducer" ;
        angle_offset_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
        angle_offset_athwartship:obligation = "NA" ;
        angle_offset_athwartship:echopype_mods = "added" ;
      double angle_sensitivity_alongship(channel, ping_time, beam) ;
        angle_sensitivity_alongship:_FillValue = NaN ;
        angle_sensitivity_alongship:long_name = "alongship angle sensitivity of the transducer" ;
        angle_sensitivity_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
        angle_sensitivity_alongship:obligation = "NA" ;
        angle_sensitivity_alongship:echopype_mods = "added" ;
      double angle_sensitivity_athwartship(channel, ping_time, beam) ;
        angle_sensitivity_athwartship:_FillValue = NaN ;
        angle_sensitivity_athwartship:long_name = "athwartship angle sensitivity of the transducer" ;
        angle_sensitivity_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
        angle_sensitivity_athwartship:obligation = "NA" ;
        angle_sensitivity_athwartship:echopype_mods = "added" ;
      float backscatter_i(channel, ping_time, range_sample, beam) ;
        backscatter_i:_FillValue = NaNf ;
        backscatter_i:long_name = "Raw backscatter measurements (imaginary part)" ;
        backscatter_i:units = "dB" ;
        backscatter_i:obligation = "MA" ;
      float backscatter_r(channel, ping_time, range_sample, beam) ;
        backscatter_r:_FillValue = NaNf ;
        backscatter_r:long_name = "Raw backscatter measurements (real part)" ;
        backscatter_r:units = "dB" ;
        backscatter_r:obligation = "M" ;
      string beam(beam) ;
        beam:long_name = "Beam name" ;
        beam:obligation = "M" ;
      double beam_direction_x(channel, ping_time, beam) ;
        beam_direction_x:_FillValue = NaN ;
        beam_direction_x:long_name = "x-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_x:units = "1" ;
        beam_direction_x:valid_range = -1., 1. ;
        beam_direction_x:obligation = "M" ;
      double beam_direction_y(channel, ping_time, beam) ;
        beam_direction_y:_FillValue = NaN ;
        beam_direction_y:long_name = "y-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_y:units = "1" ;
        beam_direction_y:valid_range = -1., 1. ;
        beam_direction_y:obligation = "M" ;
      double beam_direction_z(channel, ping_time, beam) ;
        beam_direction_z:_FillValue = NaN ;
        beam_direction_z:long_name = "z-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_z:units = "1" ;
        beam_direction_z:valid_range = -1., 1. ;
        beam_direction_z:obligation = "M" ;
      int64 beam_type(channel, ping_time) ;
        beam_type:echopype_mods = "changed-type";
        beam_type:obligation = "M" ;
      double beamwidth_twoway_alongship(channel, ping_time, beam) ;
        beamwidth_twoway_alongship:_FillValue = NaN ;
        beamwidth_twoway_alongship:long_name = "Half power two-way beam width along alongship axis of beam" ;
        beamwidth_twoway_alongship:units = "arc_degree" ;
        beamwidth_twoway_alongship:valid_range = 0., 360. ;
        beamwidth_twoway_alongship:comment = "Introduced in echopype for Simrad echosounders to avoid potential confusion with convention definitions. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. The convention defines one-way transmit or receive beamwidth (beamwidth_receive_minor and beamwidth_transmit_minor), but Simrad echosounders record two-way beamwidth in the data." ;
        beamwidth_twoway_alongship:obligation = "NA" ;
        beamwidth_twoway_alongship:echopype_mods = "added-replacement" ;
      double beamwidth_twoway_athwartship(channel, ping_time, beam) ;
        beamwidth_twoway_athwartship:_FillValue = NaN ;
        beamwidth_twoway_athwartship:long_name = "Half power two-way beam width along athwartship axis of beam" ;
        beamwidth_twoway_athwartship:units = "arc_degree" ;
        beamwidth_twoway_athwartship:valid_range = 0., 360. ;
        beamwidth_twoway_athwartship:comment = "Introduced in echopype for Simrad echosounders to avoid potential confusion with convention definitions. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. The convention defines one-way transmit or receive beamwidth (beamwidth_receive_major and beamwidth_transmit_major), but Simrad echosounders record two-way beamwidth in the data." ;
        beamwidth_twoway_athwartship:obligation = "NA" ;
        beamwidth_twoway_athwartship:echopype_mods = "added-replacement" ;
      string channel(channel) ;
        channel:long_name = "Vendor channel ID" ;
        channel:obligation = "NA" ;
        channel:echopype_mods = "added" ;
      double equivalent_beam_angle(channel, ping_time, beam) ;
        equivalent_beam_angle:_FillValue = NaN ;
        equivalent_beam_angle:long_name = "Equivalent beam angle" ;
        equivalent_beam_angle:units = "sr" ;
        equivalent_beam_angle:valid_range = 0., 12.6 ;
        equivalent_beam_angle:obligation = "M" ;
      int64 frequency_end(channel, ping_time, beam) ;
        // is this a direct replacement of transmit_frequency_end?
        frequency_end:long_name = "Ending frequency of the transducer" ;
        frequency_end:units = "Hz" ;
        frequency_end:valid_min = 0. ;
        frequency_end:standard_name = "sound_frequency" ;
        frequency_end:obligation = "NA" ;
        frequency_end:echopype_mods = "added-replacement" ;
      double frequency_nominal(channel) ;
        frequency_nominal:_FillValue = NaN ;
        frequency_nominal:units = "Hz" ;
        frequency_nominal:long_name = "Transducer frequency" ;
        frequency_nominal:valid_min = 0. ;
        frequency_nominal:standard_name = "sound_frequency" ;
        frequency_nominal:obligation = "NA" ;
        frequency_nominal:echopype_mods = "added" ;
      int64 frequency_start(channel, ping_time, beam) ;
        // is this a direct replacement of transmit_frequency_start?
        frequency_start:long_name = "Starting frequency of the transducer" ;
        frequency_start:units = "Hz" ;
        frequency_start:valid_min = 0. ;
        frequency_start:standard_name = "sound_frequency" ;
        frequency_start:obligation = "NA" ;
        frequency_start:echopype_mods = "added-replacement" ;
      double ping_time(ping_time) ;
        ping_time:_FillValue = NaN ;
        ping_time:long_name = "Timestamp of each ping" ;
        ping_time:standard_name = "time" ;
        ping_time:axis = "T" ;
        ping_time:units = "seconds since 1900-01-01T00:00:00+00:00" ;
        ping_time:calendar = "gregorian" ;
        ping_time:obligation = "M" ;
        ping_time:echopype_mods = "changed" ;
      int64 range_sample(range_sample) ;
        range_sample:long_name = "Along-range sample number, base 0" ;
        range_sample:obligation = "NA" ;
        range_sample:echopype_mods = "added" ;
      double sample_interval(channel, ping_time) ;
        sample_interval:_FillValue = NaN ;
        sample_interval:long_name = "Interval between recorded raw data samples" ;
        sample_interval:units = "s" ;
        sample_interval:valid_min = 0. ;
        sample_interval:obligation = "M" ;
      double slope(channel, ping_time) ;
        slope:_FillValue = NaN ;
        slope:echopype_mods = "added" ;
        :obligation = "M" ;
      string transceiver_software_version(channel) ;
        transceiver_software_version:obligation = "NA" ;
        transceiver_software_version:echopype_mods = "added" ;
      double transmit_power(channel, ping_time) ;
        transmit_power:_FillValue = NaN ;
        transmit_power:long_name = "Nominal transmit power" ;
        transmit_power:units = "W" ;
        transmit_power:valid_min = 0. ;
        transmit_power:obligation = "MA" ;
      float transmit_duration_nominal(channel, ping_time) ;
        transmit_duration_nominal:_FillValue = NaNf ;
        // long_name is supposed to be "Nominal duration of transmitted pulse"
        transmit_duration_nominal:long_name = "Nominal bandwidth of transmitted pulse" ;
        transmit_duration_nominal:units = "s" ;
        transmit_duration_nominal:valid_min = 0. ;
        transmit_duration_nominal:obligation = "M" ;

    // group attributes:
        :beam_mode = "vertical" ;
        :conversion_equation_t = "type_3" ;
    data:

     // --------------------------------

     angle_athwartship =
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.;

     angle_alongship =
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.,
  1., 2., 3., 4.;

     // --------------------------------

     frequency_nominal = 120000 ;

     beam_type =
  1, 1, 1, 1, 1 ;

     beamwidth_twoway_alongship =
  6.72, 6.72, 6.72, 6.72,
  6.72, 6.72, 6.72, 6.72,
  6.72, 6.72, 6.72, 6.72,
  6.72, 6.72, 6.72, 6.72,
  6.72, 6.72, 6.72, 6.72 ;

     beamwidth_twoway_athwartship =
  6.62, 6.62, 6.62, 6.62,
  6.62, 6.62, 6.62, 6.62,
  6.62, 6.62, 6.62, 6.62,
  6.62, 6.62, 6.62, 6.62,
  6.62, 6.62, 6.62, 6.62 ;

     beam_direction_x =
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;

     beam_direction_y =
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;

     beam_direction_z =
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;

     angle_offset_alongship =
  0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03 ;

     angle_offset_athwartship =
  -0.04, -0.04, -0.04, -0.04,
  -0.04, -0.04, -0.04, -0.04,
  -0.04, -0.04, -0.04, -0.04,
  -0.04, -0.04, -0.04, -0.04,
  -0.04, -0.04, -0.04, -0.04 ;

     angle_sensitivity_alongship =
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23 ;

     angle_sensitivity_athwartship =
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23,
  23, 23, 23, 23 ;

     equivalent_beam_angle =
  -20.7, -20.7, -20.7, -20.7,
  -20.7, -20.7, -20.7, -20.7,
  -20.7, -20.7, -20.7, -20.7,
  -20.7, -20.7, -20.7, -20.7,
  -20.7, -20.7, -20.7, -20.7 ;

     transceiver_software_version = "2.20" ;

     channel = "WBT 150013-15 ES120-7C_ES" ;

     backscatter_r =
  3.748114e-05, 3.223628e-05, 4.797172e-05, 4.606434e-05,
  -0.001821251, -0.001401654, -0.002360794, -0.002269238,
  -0.004355508, -0.004630208, -0.004447064, -0.005667772,
  9.937377e-06, -0.002696561, 0.001752623, -0.001180428,
  0.001786956, 0.001405496, 0.0002138335, 0.0009125524,
  -0.001535143, -0.0003694827, -0.001317735, -0.0008839236,
  0.0008839405, -0.0002760307, 0.005576149, 0.001294855,
  -0.004096094, -0.0004257597, -0.008436286, -0.005194717,
  -0.004813255, -0.002467665, -0.003657839, 0.0003294374,
  0.005087816, 0.002383663, 0.009992199, 0.008527683;
  
     backscatter_i =
  -1.39895e-05, -2.619089e-05, 9.81713e-06, -8.684628e-06,
  -0.001550432, -0.0006722168, -0.002749895, -0.002154805,
  -0.006812171, -0.002261649, -0.01240351, -0.008802476,
  -0.005438801, -0.00137876, -0.00895407, -0.00565234,
  0.004050044, 0.002032642, 0.006811983, 0.005804872,
  -0.0004639029, -0.001512256, -0.002994009, -0.002627701,
  -0.002833841, -0.001790773, -0.004935201, -0.004935273,
  0.005743994, 0.005377867, 0.008619457, 0.00819222,
  0.0006874841, 0.001214742, -0.0007828317, 0.001909023,
  0.007132462, 0.005392954, 0.008863428, 0.006247404;
  

     ping_time = 3842381772.962, 3842381773.963, 3842381774.965, 
        3842381775.962, 3842381776.964 ;

     range_sample = 0, 1 ;

     beam = "1", "2", "3", "4" ;

     frequency_start =
  90000, 90000, 90000, 90000,
  90000, 90000, 90000, 90000,
  90000, 90000, 90000, 90000,
  90000, 90000, 90000, 90000,
  90000, 90000, 90000, 90000 ;

     frequency_end =
  170000, 170000, 170000, 170000,
  170000, 170000, 170000, 170000,
  170000, 170000, 170000, 170000,
  170000, 170000, 170000, 170000,
  170000, 170000, 170000, 170000 ;

     sample_interval =
  8e-06, 8e-06, 8e-06, 8e-06, 8e-06 ;

     transmit_power =
  50, 50, 50, 50, 50 ;

     transmit_duration_nominal =
  0.000512, 0.000512, 0.000512, 0.000512, 0.000512 ;

     slope =
  0.5, 0.5, 0.5, 0.5, 0.5 ;
    } // group Beam_group1

  group: Beam_group2 {
    dimensions:
      channel = 2 ;
      ping_time = 5 ;
      beam = 1 ;
      range_sample = 2 ;
    variables:
      double frequency_nominal(channel) ;
        frequency_nominal:_FillValue = NaN ;
        frequency_nominal:units = "Hz" ;
        frequency_nominal:long_name = "Transducer frequency" ;
        frequency_nominal:valid_min = 0. ;
        frequency_nominal:standard_name = "sound_frequency" ;
      int64 beam_type(channel, ping_time) ;
      double beamwidth_twoway_alongship(channel, ping_time, beam) ;
        beamwidth_twoway_alongship:_FillValue = NaN ;
        beamwidth_twoway_alongship:long_name = "Half power two-way beam width along alongship axis of beam" ;
        beamwidth_twoway_alongship:units = "arc_degree" ;
        beamwidth_twoway_alongship:valid_range = 0., 360. ;
        beamwidth_twoway_alongship:comment = "Introduced in echopype for Simrad echosounders to avoid potential confusion with convention definitions. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. The convention defines one-way transmit or receive beamwidth (beamwidth_receive_minor and beamwidth_transmit_minor), but Simrad echosounders record two-way beamwidth in the data." ;
      double beamwidth_twoway_athwartship(channel, ping_time, beam) ;
        beamwidth_twoway_athwartship:_FillValue = NaN ;
        beamwidth_twoway_athwartship:long_name = "Half power two-way beam width along athwartship axis of beam" ;
        beamwidth_twoway_athwartship:units = "arc_degree" ;
        beamwidth_twoway_athwartship:valid_range = 0., 360. ;
        beamwidth_twoway_athwartship:comment = "Introduced in echopype for Simrad echosounders to avoid potential confusion with convention definitions. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. The convention defines one-way transmit or receive beamwidth (beamwidth_receive_major and beamwidth_transmit_major), but Simrad echosounders record two-way beamwidth in the data." ;
      double beam_direction_x(channel, ping_time, beam) ;
        beam_direction_x:_FillValue = NaN ;
        beam_direction_x:long_name = "x-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_x:units = "1" ;
        beam_direction_x:valid_range = -1., 1. ;
      double beam_direction_y(channel, ping_time, beam) ;
        beam_direction_y:_FillValue = NaN ;
        beam_direction_y:long_name = "y-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_y:units = "1" ;
        beam_direction_y:valid_range = -1., 1. ;
      double beam_direction_z(channel, ping_time, beam) ;
        beam_direction_z:_FillValue = NaN ;
        beam_direction_z:long_name = "z-component of the vector that gives the pointing direction of the beam, in sonar beam coordinate system" ;
        beam_direction_z:units = "1" ;
        beam_direction_z:valid_range = -1., 1. ;
      double angle_offset_alongship(channel, ping_time, beam) ;
        angle_offset_alongship:_FillValue = NaN ;
        angle_offset_alongship:long_name = "electrical alongship angle offset of the transducer" ;
        angle_offset_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
      double angle_offset_athwartship(channel, ping_time, beam) ;
        angle_offset_athwartship:_FillValue = NaN ;
        angle_offset_athwartship:long_name = "electrical athwartship angle offset of the transducer" ;
        angle_offset_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
      double angle_sensitivity_alongship(channel, ping_time, beam) ;
        angle_sensitivity_alongship:_FillValue = NaN ;
        angle_sensitivity_alongship:long_name = "alongship angle sensitivity of the transducer" ;
        angle_sensitivity_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
      double angle_sensitivity_athwartship(channel, ping_time, beam) ;
        angle_sensitivity_athwartship:_FillValue = NaN ;
        angle_sensitivity_athwartship:long_name = "athwartship angle sensitivity of the transducer" ;
        angle_sensitivity_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
      double equivalent_beam_angle(channel, ping_time, beam) ;
        equivalent_beam_angle:_FillValue = NaN ;
        equivalent_beam_angle:long_name = "Equivalent beam angle" ;
        equivalent_beam_angle:units = "sr" ;
        equivalent_beam_angle:valid_range = 0., 12.5663706143592 ;
      string transceiver_software_version(channel) ;
      string channel(channel) ;
        channel:long_name = "Vendor channel ID" ;
      float backscatter_r(channel, ping_time, range_sample, beam) ;
        backscatter_r:_FillValue = NaNf ;
        backscatter_r:long_name = "Backscatter power" ;
        backscatter_r:units = "dB" ;
      double ping_time(ping_time) ;
        ping_time:_FillValue = NaN ;
        ping_time:long_name = "Timestamp of each ping" ;
        ping_time:standard_name = "time" ;
        ping_time:axis = "T" ;
        ping_time:units = "seconds since 1900-01-01T00:00:00+00:00" ;
        ping_time:calendar = "gregorian" ;
      int64 range_sample(range_sample) ;
        range_sample:long_name = "Along-range sample number, base 0" ;
      double angle_athwartship(channel, ping_time, range_sample, beam) ;
        angle_athwartship:_FillValue = NaN ;
        angle_athwartship:long_name = "electrical athwartship angle" ;
        angle_athwartship:comment = "Introduced in echopype for Simrad echosounders. The athwartship angle corresponds to the major angle in SONAR-netCDF4 vers 2. " ;
      double angle_alongship(channel, ping_time, range_sample, beam) ;
        angle_alongship:_FillValue = NaN ;
        angle_alongship:long_name = "electrical alongship angle" ;
        angle_alongship:comment = "Introduced in echopype for Simrad echosounders. The alongship angle corresponds to the minor angle in SONAR-netCDF4 vers 2. " ;
      double sample_interval(channel, ping_time) ;
        sample_interval:_FillValue = NaN ;
        sample_interval:long_name = "Interval between recorded raw data samples" ;
        sample_interval:units = "s" ;
        sample_interval:valid_min = 0. ;
      double transmit_power(channel, ping_time) ;
        transmit_power:_FillValue = NaN ;
        transmit_power:long_name = "Nominal transmit power" ;
        transmit_power:units = "W" ;
        transmit_power:valid_min = 0. ;
      float transmit_duration_nominal(channel, ping_time) ;
        transmit_duration_nominal:_FillValue = NaNf ;
        transmit_duration_nominal:long_name = "Nominal bandwidth of transmitted pulse" ;
        transmit_duration_nominal:units = "s" ;
        transmit_duration_nominal:valid_min = 0. ;
      double slope(channel, ping_time) ;
        slope:_FillValue = NaN ;
      string beam(beam) ;
        beam:long_name = "Beam name" ;

    // group attributes:
        :beam_mode = "vertical" ;
        :conversion_equation_t = "type_3" ;
    data:

     frequency_nominal = 200000, 70000 ;

     beam_type =
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1 ;

     beamwidth_twoway_alongship =
  7.47,
  7.47,
  7.47,
  7.47,
  7.47,
  6.86,
  6.86,
  6.86,
  6.86,
  6.86 ;

     beamwidth_twoway_athwartship =
  6.9,
  6.9,
  6.9,
  6.9,
  6.9,
  6.65,
  6.65,
  6.65,
  6.65,
  6.65 ;

     beam_direction_x =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

     beam_direction_y =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

     beam_direction_z =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

     angle_offset_alongship =
  -0.14,
  -0.14,
  -0.14,
  -0.14,
  -0.14,
  0.03,
  0.03,
  0.03,
  0.03,
  0.03 ;

     angle_offset_athwartship =
  -0.17,
  -0.17,
  -0.17,
  -0.17,
  -0.17,
  0.06,
  0.06,
  0.06,
  0.06,
  0.06 ;

     angle_sensitivity_alongship =
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23 ;

     angle_sensitivity_athwartship =
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23,
  23 ;

     equivalent_beam_angle =
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7,
  -20.7 ;

     transceiver_software_version = "2.20", "2.20" ;

     channel = "WBT 545612-15 ES200-7C_ES", "WBT 549762-15 ES70-7C_ES" ;

     backscatter_r =
  -37.86393,
  -53.9267,
  -62.82825,
  -64.34516,
  -54.90269,
  -89.6505,
  -147.9515,
  -151.7027,
  -148.1279,
  -156.2416,
  -152.173,
  -136.2631,
  -138.2621,
  -154.3719,
  -150.7972,
  -143.7418,
  -137.1685,
  -126.6795,
  -127.5732,
  -146.5052 ;

     ping_time = 3842381772.962, 3842381773.963, 3842381774.965, 
        3842381775.962, 3842381776.964 ;

     range_sample = 0, 1 ;

     angle_athwartship =
  -8,
  111,
  112,
  -108,
  48,
  61,
  54,
  -39,
  -2,
  -52,
  11,
  28,
  47,
  -65,
  -104,
  -5,
  93,
  -28,
  114,
  124 ;

     angle_alongship =
  0,
  -78,
  93,
  70,
  54,
  -102,
  27,
  -33,
  -46,
  -99,
  -127,
  67,
  -7,
  -116,
  -124,
  -8,
  -14,
  -7,
  -120,
  109 ;

     sample_interval =
  0.00012, 0.00012, 0.00012, 0.00012, 0.00012,
  0.00012, 0.00012, 0.00012, 0.00012, 0.00012 ;

     transmit_power =
  45, 45, 45, 45, 45,
  75, 75, 75, 75, 75 ;

     transmit_duration_nominal =
  0.000512, 0.000512, 0.000512, 0.000512, 0.000512,
  0.000512, 0.000512, 0.000512, 0.000512, 0.000512 ;

     slope =
  0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5 ;

     beam = "1" ;
    } // group Beam_group2
  } // group Sonar

group: Vendor_specific {
  dimensions:
    channel = 3 ;
    pulse_length_bin = 5 ;
  variables:
    double frequency_nominal(channel) ;
      frequency_nominal:_FillValue = NaN ;
      frequency_nominal:units = "Hz" ;
      frequency_nominal:long_name = "Transducer frequency" ;
      frequency_nominal:valid_min = 0. ;
      frequency_nominal:standard_name = "sound_frequency" ;
    double sa_correction(channel, pulse_length_bin) ;
      sa_correction:_FillValue = NaN ;
    double gain_correction(channel, pulse_length_bin) ;
      gain_correction:_FillValue = NaN ;
    double pulse_length(channel, pulse_length_bin) ;
      pulse_length:_FillValue = NaN ;
    string channel(channel) ;
      channel:long_name = "Vendor channel ID" ;
    int64 pulse_length_bin(pulse_length_bin) ;
    int64 impedance_transceiver(channel) ;
      impedance_transceiver:units = "ohm" ;
      impedance_transceiver:long_name = "Transceiver impedance" ;
    double fs_receiver(channel) ;
      fs_receiver:_FillValue = NaN ;
      fs_receiver:units = "Hz" ;
      fs_receiver:long_name = "Receiver sampling frequency" ;
    string transceiver_type(channel) ;
      transceiver_type:long_name = "Transceiver type" ;

  // group attributes:
      :WBT\ 150013-15\ ES120-7C_ES\ WBT\ filter_r = 6.497843e-05f, 0.0004637341f, 0.0006013685f, -0.001046955f, -0.006130705f, -0.01373757f, -0.01884355f, -0.01544923f, -0.004006708f, 0.003928663f, -0.007787384f, -0.04297968f, -0.07997828f, -0.07907871f, -0.01193036f, 0.1085594f, 0.2261203f, 0.2749873f, 0.2261203f, 0.1085594f, -0.01193036f, -0.07907871f, -0.07997828f, -0.04297968f, -0.007787384f, 0.003928663f, -0.004006708f, -0.01544923f, -0.01884355f, -0.01373757f, -0.006130705f, -0.001046955f, 0.0006013685f, 0.0004637341f, 6.497843e-05f ;
      :WBT\ 150013-15\ ES120-7C_ES\ WBT\ filter_i = 1.099028e-05f, 0.0004002846f, 0.001850822f, 0.004463713f, 0.00626047f, 0.003527209f, -0.005689203f, -0.01715811f, -0.0210039f, -0.01056386f, 0.006172204f, 0.005429597f, -0.03560863f, -0.1137794f, -0.1896276f, -0.207655f, -0.1369433f, 0.f, 0.1369433f, 0.207655f, 0.1896276f, 0.1137794f, 0.03560863f, -0.005429597f, -0.006172204f, 0.01056386f, 0.0210039f, 0.01715811f, 0.005689203f, -0.003527209f, -0.00626047f, -0.004463713f, -0.001850822f, -0.0004002846f, -1.099028e-05f ;
      :WBT\ 150013-15\ ES120-7C_ES\ PC\ filter_r = 4.295626e-05f, -0.0002459195f, 0.0006159935f, -0.0009566006f, 0.0008330459f, -0.0001137168f, -0.0007683993f, 0.0009682976f, -0.0001464992f, -0.001003838f, 0.001241533f, -0.0001291441f, -0.001300661f, 0.001486752f, -8.421461e-05f, -0.001489456f, 0.001539964f, -1.387342e-05f, -0.001403014f, 0.001252724f, 4.82855e-05f, -0.0008746417f, 0.000529956f, 2.176987e-05f, 0.0002278514f, -0.0006306252f, -0.0002104291f, 0.001952389f, -0.002115786f, -0.0007595157f, 0.004200612f, -0.00368967f, -0.001677608f, 0.006688344f, -0.005024858f, -0.002894634f, 0.008938159f, -0.005769955f, -0.004157946f, 0.01030561f, -0.005632245f, -0.004998442f, 0.01004108f, -0.004463988f, -0.00471662f, 0.007351779f, -0.002326037f, -0.002356081f, 0.00138546f, 0.0005019079f, 0.003439446f, -0.009041226f, 0.003558592f, 0.01514272f, -0.02672362f, 0.006292708f, 0.04008081f, -0.06336121f, 0.00818312f, 0.1287748f, -0.2777138f, 0.3422951f, -0.2777138f, 0.1287748f, 0.00818312f, -0.06336121f, 0.04008081f, 0.006292708f, -0.02672362f, 0.01514272f, 0.003558592f, -0.009041226f, 0.003439447f, 0.0005019079f, 0.00138546f, -0.002356081f, -0.002326037f, 0.007351779f, -0.00471662f, -0.004463988f, 0.01004108f, -0.004998442f, -0.005632245f, 0.01030561f, -0.004157946f, -0.005769955f, 0.008938159f, -0.002894634f, -0.005024858f, 0.006688344f, -0.001677608f, -0.00368967f, 0.004200612f, -0.0007595157f, -0.002115786f, 0.001952389f, -0.0002104291f, -0.0006306252f, 0.0002278514f, 2.176987e-05f, 0.000529956f, -0.0008746417f, 4.82855e-05f, 0.001252724f, -0.001403014f, -1.387342e-05f, 0.001539964f, -0.001489456f, -8.421461e-05f, 0.001486752f, -0.001300661f, -0.0001291441f, 0.001241533f, -0.001003838f, -0.0001464992f, 0.0009682976f, -0.0007683993f, -0.0001137168f, 0.0008330459f, -0.0009566006f, 0.0006159935f, -0.0002459195f, 4.295626e-05f ;
      :WBT\ 150013-15\ ES120-7C_ES\ PC\ filter_i = -0.0002223318f, 0.0007585372f, -0.001307896f, 0.001508219f, -0.001006322f, 0.0001072982f, 0.0005586701f, -0.0005320269f, 5.821858e-05f, 0.0002578815f, -0.0001567734f, 1.240506e-13f, -0.0001643805f, 0.0003815934f, -3.355839e-05f, -0.0008191344f, 0.001118454f, -1.353905e-05f, -0.00169661f, 0.001973119f, 0.0001014554f, -0.002693545f, 0.002775274f, 0.0003373723f, -0.003612944f, 0.003308706f, 0.0006493092f, -0.004147882f, 0.003334803f, 0.0009187546f, -0.003944126f, 0.002681097f, 0.0009225718f, -0.002647887f, 0.001290304f, 0.0003657461f, -8.585729e-12f, -0.0007289836f, -0.001067719f, 0.004080063f, -0.003096652f, -0.003631976f, 0.009428687f, -0.005396692f, -0.007433061f, 0.01562217f, -0.007160481f, -0.01235386f, 0.02201261f, -0.007968948f, -0.01802736f, 0.02782771f, -0.007561236f, -0.02386025f, 0.03230396f, -0.005908735f, -0.02912002f, 0.03483342f, -0.003239711f, -0.03306362f, 0.03508348f, -3.28802e-10f, -0.03508348f, 0.03306362f, 0.003239711f, -0.03483342f, 0.02912002f, 0.005908735f, -0.03230396f, 0.02386025f, 0.007561236f, -0.02782771f, 0.01802736f, 0.007968948f, -0.02201261f, 0.01235386f, 0.007160481f, -0.01562217f, 0.007433061f, 0.005396692f, -0.009428687f, 0.003631976f, 0.003096652f, -0.004080063f, 0.001067719f, 0.0007289837f, -8.585913e-12f, -0.0003657461f, -0.001290304f, 0.002647887f, -0.0009225718f, -0.002681097f, 0.003944126f, -0.0009187546f, -0.003334803f, 0.004147882f, -0.0006493092f, -0.003308706f, 0.003612944f, -0.0003373723f, -0.002775274f, 0.002693545f, -0.0001014554f, -0.001973119f, 0.00169661f, 1.353905e-05f, -0.001118454f, 0.0008191344f, 3.355839e-05f, -0.0003815934f, 0.0001643805f, 1.240559e-13f, 0.0001567734f, -0.0002578815f, -5.821858e-05f, 0.0005320269f, -0.0005586701f, -0.0001072982f, 0.001006322f, -0.001508219f, 0.001307896f, -0.0007585372f, 0.0002223318f ;
      :WBT\ 545612-15\ ES200-7C_ES\ WBT\ filter_r = 0.0001670101f, 0.0003854856f, 0.0002711259f, -0.0008084571f, -0.002679517f, -0.003521757f, -0.0006867192f, 0.006353701f, 0.01322204f, 0.01192107f, -0.002436285f, -0.02401397f, -0.03607074f, -0.02238351f, 0.01643263f, 0.05652861f, 0.06449548f, 0.02442409f, -0.04343958f, -0.09176075f, -0.08053276f, -0.01085334f, 0.07125145f, 0.1073812f, 0.07125145f, -0.01085334f, -0.08053276f, -0.09176075f, -0.04343958f, 0.02442409f, 0.06449548f, 0.05652861f, 0.01643263f, -0.02238351f, -0.03607074f, -0.02401397f, -0.002436285f, 0.01192107f, 0.01322204f, 0.006353701f, -0.0006867192f, -0.003521757f, -0.002679517f, -0.0008084571f, 0.0002711259f, 0.0003854856f, 0.0001670101f ;
      :WBT\ 545612-15\ ES200-7C_ES\ WBT\ filter_i = -7.43577e-05f, 0.0001716292f, 0.0008344396f, 0.001400289f, 0.0005695489f, -0.002558706f, -0.006533697f, -0.007056499f, 6.47693e-18f, 0.01323969f, 0.0231797f, 0.01744717f, -0.007667072f, -0.03876937f, -0.05057442f, -0.02516816f, 0.02871524f, 0.07516961f, 0.07523956f, 0.01950435f, -0.05851047f, -0.1032627f, -0.07913276f, 0.f, 0.07913276f, 0.1032627f, 0.05851047f, -0.01950435f, -0.07523956f, -0.07516961f, -0.02871524f, 0.02516816f, 0.05057442f, 0.03876937f, 0.007667072f, -0.01744717f, -0.0231797f, -0.01323969f, -6.47693e-18f, 0.007056499f, 0.006533697f, 0.002558706f, -0.0005695489f, -0.001400289f, -0.0008344396f, -0.0001716292f, 7.43577e-05f ;
      :WBT\ 545612-15\ ES200-7C_ES\ PC\ filter_r = -4.927609e-05f, 3.760648e-05f, 0.0002431257f, 0.0001341616f, -0.0005857545f, -0.000920431f, 0.000527535f, 0.002469935f, 0.001067847f, -0.003802111f, -0.005036109f, 0.002488046f, 0.0101937f, 0.003907911f, -0.01245748f, -0.01489876f, 0.006691383f, 0.02505566f, 0.00882041f, -0.02591737f, -0.02866697f, 0.01194079f, 0.04156194f, 0.01362727f, -0.03735335f, -0.03859383f, 0.0150322f, 0.04896387f, 0.0150322f, -0.03859383f, -0.03735336f, 0.01362727f, 0.04156194f, 0.01194079f, -0.02866697f, -0.02591737f, 0.00882041f, 0.02505566f, 0.006691383f, -0.01489876f, -0.01245748f, 0.003907911f, 0.0101937f, 0.002488046f, -0.005036109f, -0.003802111f, 0.001067847f, 0.002469935f, 0.0005275351f, -0.000920431f, -0.0005857545f, 0.0001341616f, 0.0002431257f, 3.760648e-05f, -4.927609e-05f ;
      :WBT\ 545612-15\ ES200-7C_ES\ PC\ filter_i = 3.553911e-05f, 0.000116851f, 1.770665e-12f, -0.000414017f, -0.0004253135f, 0.0006684702f, 0.001624696f, 1.798833e-11f, -0.003287604f, -0.002762133f, 0.003658685f, 0.007658527f, 7.423982e-11f, -0.01202842f, -0.009050624f, 0.01082432f, 0.02059507f, 1.82478e-10f, -0.02714754f, -0.01882981f, 0.02082751f, 0.03675107f, 3.026916e-10f, -0.04194153f, -0.02713854f, 0.0280398f, 0.04626546f, 3.565989e-10f, -0.04626546f, -0.0280398f, 0.02713854f, 0.04194153f, 3.026912e-10f, -0.03675107f, -0.02082751f, 0.01882981f, 0.02714754f, 1.824776e-10f, -0.02059507f, -0.01082432f, 0.009050624f, 0.01202842f, 7.423948e-11f, -0.007658527f, -0.003658685f, 0.002762133f, 0.003287604f, 1.798824e-11f, -0.001624696f, -0.0006684702f, 0.0004253135f, 0.000414017f, 1.770656e-12f, -0.000116851f, -3.553911e-05f ;
      :WBT\ 549762-15\ ES70-7C_ES\ WBT\ filter_r = 0.0001637498f, 0.0004160573f, 0.0008704634f, 0.001477125f, 0.002073696f, 0.002332524f, 0.001766719f, -0.0001988578f, -0.004085834f, -0.0101677f, -0.01826584f, -0.02759846f, -0.03674725f, -0.04378875f, -0.04659944f, -0.04329395f, -0.03270828f, -0.01481024f, 0.009081345f, 0.03635313f, 0.06345171f, 0.08648343f, 0.1019389f, 0.1073812f, 0.1019389f, 0.08648343f, 0.06345171f, 0.03635313f, 0.009081345f, -0.01481024f, -0.03270828f, -0.04329395f, -0.04659944f, -0.04378875f, -0.03674725f, -0.02759846f, -0.01826584f, -0.0101677f, -0.004085834f, -0.0001988578f, 0.001766719f, 0.002332524f, 0.002073696f, 0.001477125f, 0.0008704634f, 0.0004160573f, 0.0001637498f ;
      :WBT\ 549762-15\ ES70-7C_ES\ WBT\ filter_i = -8.128613e-05f, -7.037082e-05f, 0.0001099651f, 0.0006576583f, 0.001789967f, 0.00367547f, 0.006327676f, 0.009493374f, 0.0125749f, 0.0146294f, 0.01447733f, 0.010927f, 0.003085753f, -0.009307585f, -0.02561826f, -0.04421033f, -0.06256517f, -0.07763802f, -0.08640323f, -0.08648067f, -0.07669994f, -0.05745946f, -0.03077715f, 0.f, 0.03077715f, 0.05745946f, 0.07669994f, 0.08648067f, 0.08640323f, 0.07763802f, 0.06256517f, 0.04421033f, 0.02561826f, 0.009307585f, -0.003085753f, -0.010927f, -0.01447733f, -0.0146294f, -0.0125749f, -0.009493374f, -0.006327676f, -0.00367547f, -0.001789967f, -0.0006576583f, -0.0001099651f, 7.037082e-05f, 8.128613e-05f ;
      :WBT\ 549762-15\ ES70-7C_ES\ PC\ filter_r = -5.551979e-05f, -2.232542e-05f, 0.0002441836f, -8.08744e-05f, -0.000672077f, 0.0006100768f, 0.001246f, -0.001997815f, -0.001471134f, 0.004552286f, 0.0003915385f, -0.007988461f, 0.003150835f, 0.01108373f, -0.009814262f, -0.01173775f, 0.01897707f, 0.007743436f, -0.02831885f, 0.002012204f, 0.03432137f, -0.01645243f, -0.03362393f, 0.03214819f, 0.02474028f, -0.04435353f, -0.009114732f, 0.04896496f, -0.009114732f, -0.04435353f, 0.02474028f, 0.03214819f, -0.03362393f, -0.01645243f, 0.03432137f, 0.002012204f, -0.02831885f, 0.007743436f, 0.01897707f, -0.01173775f, -0.009814262f, 0.01108373f, 0.003150835f, -0.007988461f, 0.0003915386f, 0.004552286f, -0.001471134f, -0.001997815f, 0.001246f, 0.0006100768f, -0.000672077f, -8.087439e-05f, 0.0002441836f, -2.232542e-05f, -5.551979e-05f ;
      :WBT\ 549762-15\ ES70-7C_ES\ PC\ filter_i = 2.225783e-05f, -0.0001206882f, 7.97766e-13f, 0.0004276127f, -0.0002663701f, -0.0009602288f, 0.001169417f, 0.001452004f, -0.0031278f, -0.001168649f, 0.006212248f, -0.001009265f, -0.009695129f, 0.00609295f, 0.01186425f, -0.01418934f, -0.01043235f, 0.0238297f, 0.00357759f, -0.03197199f, 0.008812051f, 0.03496468f, -0.02442972f, -0.0301885f, 0.03898335f, 0.01756108f, -0.04778475f, 1.599717e-10f, 0.04778475f, -0.01756108f, -0.03898335f, 0.0301885f, 0.02442972f, -0.03496468f, -0.008812051f, 0.03197199f, -0.00357759f, -0.0238297f, 0.01043235f, 0.01418934f, -0.01186425f, -0.00609295f, 0.009695129f, 0.001009265f, -0.006212248f, 0.001168649f, 0.0031278f, -0.001452004f, -0.001169417f, 0.0009602288f, 0.0002663701f, -0.0004276127f, 7.977617e-13f, 0.0001206882f, -2.225783e-05f ;
      :WBT\ 150013-15\ ES120-7C_ES\ WBT\ decimation = 6LL ;
      :WBT\ 150013-15\ ES120-7C_ES\ PC\ decimation = 2LL ;
      :WBT\ 545612-15\ ES200-7C_ES\ WBT\ decimation = 6LL ;
      :WBT\ 545612-15\ ES200-7C_ES\ PC\ decimation = 3LL ;
      :WBT\ 549762-15\ ES70-7C_ES\ WBT\ decimation = 6LL ;
      :WBT\ 549762-15\ ES70-7C_ES\ PC\ decimation = 3LL ;
      :config_xml = "<?xml version=\"1.0\" encoding=\"utf-8\" ?>\n<Configuration>\n    <Header Copyright=\"Copyright(c) Kongsberg Maritime AS, Norway\" ApplicationName=\"EK80\" Version=\"2.0.1.0\" FileFormatVersion=\"1.23\" TimeBias=\"420\" />\n    <ActivePingMode Mode=\"Direct\" />\n    <Transceivers MergeOperation=\"AddNodeTree\">\n        <Transceiver TransceiverName=\"WBT 549762\" IPAddress=\"157.237.15.100\" MarketSegment=\"Scientific\" SerialNumber=\"549762\" Impedance=\"5400\" Multiplexing=\"0\" RxSampleFrequency=\"1500000\" EthernetAddress=\"009072086382\" Version=\"[0] Ethernet: 00:90:72:08:63:82&#x0D;&#x0A;[1] Parts-list: WBT 371790/D&#x0D;&#x0A;[2] Product: WBT&#x0D;&#x0A;IP Address: 157.237.15.100&#x0D;&#x0A;Subnet mask: 255.255.0.0&#x0D;&#x0A;Default gateway: 157.237.15.1&#x0D;&#x0A;Serial number: 549762&#x0D;&#x0A;Embedded software: Rev. 2.20&#x0D;&#x0A;FPGA TX firmware: Rev. 4&#x0D;&#x0A;FPGA RX firmware: Rev. 7&#x0D;&#x0A;CH1: 520W CH2: 508W CH3: 499W CH4: 504W&#x0D;&#x0A;TRD1: Unable to detect transducer&#x0D;&#x0A;TRD2: Unable to detect transducer&#x0D;&#x0A;TRD3: Unable to detect transducer&#x0D;&#x0A;TRD4: Unable to detect transducer&#x0D;&#x0A;\" TransceiverSoftwareVersion=\"2.20\" TransceiverNumber=\"1\" TransceiverType=\"WBT\">\n            <Channels>\n                <Channel ChannelID=\"WBT 549762-15 ES70-7C_ES\" LogicalChannelID=\"WBT 549762-15 ES70-7C\" ChannelIdShort=\"ES70-7C Serial No: 116\" MaxTxPowerTransceiver=\"2000\" HWChannelConfiguration=\"15\" PulseDuration=\"0.000128;0.000256;0.000512;0.001024;0.002048\" PulseDurationFM=\"0.000512;0.001024;0.002048;0.004096;0.008192\">\n                    <Transducer TransducerName=\"ES70-7C\" SerialNumber=\"116\" Frequency=\"70000\" FrequencyMinimum=\"45000\" FrequencyMaximum=\"90000\" MaxTxPowerTransducer=\"750\" Gain=\"27;27;27;28.88;27\" SaCorrection=\"0;0;0;-0.02;0\" EquivalentBeamAngle=\"-20.7\" DirectivityDropAt2XBeamWidth=\"0\" AngleSensitivityAlongship=\"23\" AngleSensitivityAthwartship=\"23\" AngleOffsetAlongship=\"0.03\" AngleOffsetAthwartship=\"0.06\" BeamWidthAlongship=\"6.86\" BeamWidthAthwartship=\"6.65\" BeamType=\"1\" />\n                </Channel>\n            </Channels>\n        </Transceiver>\n        <Transceiver TransceiverName=\"WBT 150013\" IPAddress=\"157.237.15.102\" MarketSegment=\"Scientific\" SerialNumber=\"150013\" Impedance=\"5400\" Multiplexing=\"0\" RxSampleFrequency=\"1500000\" EthernetAddress=\"0090720249fd\" Version=\"[0] Ethernet: 00:90:72:02:49:FD&#x0D;&#x0A;[1] Parts-list: WBT 371790/F&#x0D;&#x0A;[2] Product: WBT&#x0D;&#x0A;IP Address: 157.237.15.102&#x0D;&#x0A;Subnet mask: 255.255.0.0&#x0D;&#x0A;Default gateway: 157.237.15.1&#x0D;&#x0A;Serial number: 150013&#x0D;&#x0A;Embedded software: Rev. 2.20&#x0D;&#x0A;FPGA TX firmware: Rev. 5&#x0D;&#x0A;FPGA RX firmware: Rev. 7&#x0D;&#x0A;CH1: 502W CH2: 497W CH3: 479W CH4: 488W&#x0D;&#x0A;TRD1: Unable to detect transducer&#x0D;&#x0A;TRD2: Unable to detect transducer&#x0D;&#x0A;TRD3: Unable to detect transducer&#x0D;&#x0A;TRD4: Unable to detect transducer&#x0D;&#x0A;\" TransceiverSoftwareVersion=\"2.20\" TransceiverNumber=\"2\" TransceiverType=\"WBT\">\n            <Channels>\n                <Channel ChannelID=\"WBT 150013-15 ES120-7C_ES\" LogicalChannelID=\"WBT 150013-15 ES120-7C\" ChannelIdShort=\"ES120-7C Serial No: 1808\" MaxTxPowerTransceiver=\"2000\" HWChannelConfiguration=\"15\" PulseDuration=\"6.4e-05;0.000128;0.000256;0.000512;0.001024\" PulseDurationFM=\"0.000512;0.001024;0.002048;0.004096;0.008192\">\n                    <Transducer TransducerName=\"ES120-7C\" SerialNumber=\"1808\" Frequency=\"120000\" FrequencyMinimum=\"90000\" FrequencyMaximum=\"170000\" MaxTxPowerTransducer=\"250\" Gain=\"27;27;27;27;27.12\" SaCorrection=\"0;0;0;0;-0.08\" EquivalentBeamAngle=\"-20.7\" DirectivityDropAt2XBeamWidth=\"0\" AngleSensitivityAlongship=\"23\" AngleSensitivityAthwartship=\"23\" AngleOffsetAlongship=\"0.03\" AngleOffsetAthwartship=\"-0.04\" BeamWidthAlongship=\"6.72\" BeamWidthAthwartship=\"6.62\" BeamType=\"1\" />\n                </Channel>\n            </Channels>\n        </Transceiver>\n        <Transceiver TransceiverName=\"WBT 545612\" IPAddress=\"157.237.15.101\" MarketSegment=\"Scientific\" SerialNumber=\"545612\" Impedance=\"5400\" Multiplexing=\"0\" RxSampleFrequency=\"1500000\" EthernetAddress=\"00907208534c\" Version=\"[0] Ethernet: 00:90:72:08:53:4C&#x0D;&#x0A;[1] Parts-list: WBT 371790/D&#x0D;&#x0A;[2] Product: WBT&#x0D;&#x0A;IP Address: 157.237.15.101&#x0D;&#x0A;Subnet mask: 255.255.0.0&#x0D;&#x0A;Default gateway: 157.237.15.1&#x0D;&#x0A;Serial number: 545612&#x0D;&#x0A;Embedded software: Rev. 2.20&#x0D;&#x0A;FPGA TX firmware: Rev. 4&#x0D;&#x0A;FPGA RX firmware: Rev. 7&#x0D;&#x0A;CH1: 515W CH2: 499W CH3: 491W CH4: 499W&#x0D;&#x0A;TRD1: Unable to detect transducer&#x0D;&#x0A;TRD2: Unable to detect transducer&#x0D;&#x0A;TRD3: Unable to detect transducer&#x0D;&#x0A;TRD4: Unable to detect transducer&#x0D;&#x0A;\" TransceiverSoftwareVersion=\"2.20\" TransceiverNumber=\"3\" TransceiverType=\"WBT\">\n            <Channels>\n                <Channel ChannelID=\"WBT 545612-15 ES200-7C_ES\" LogicalChannelID=\"WBT 545612-15 ES200-7C\" ChannelIdShort=\"ES200-7C Serial No: 213\" MaxTxPowerTransceiver=\"2000\" HWChannelConfiguration=\"15\" PulseDuration=\"6.4e-05;0.000128;0.000256;0.000512;0.001024\" PulseDurationFM=\"0.000512;0.001024;0.002048;0.004096;0.008192\">\n                    <Transducer TransducerName=\"ES200-7C\" SerialNumber=\"213\" Frequency=\"200000\" FrequencyMinimum=\"160000\" FrequencyMaximum=\"260000\" MaxTxPowerTransducer=\"150\" Gain=\"26;26;26;26;26.84\" SaCorrection=\"0;0;0;0;-0.02\" EquivalentBeamAngle=\"-20.7\" DirectivityDropAt2XBeamWidth=\"0\" AngleSensitivityAlongship=\"23\" AngleSensitivityAthwartship=\"23\" AngleOffsetAlongship=\"-0.14\" AngleOffsetAthwartship=\"-0.17\" BeamWidthAlongship=\"7.47\" BeamWidthAthwartship=\"6.9\" BeamType=\"1\" />\n                </Channel>\n            </Channels>\n        </Transceiver>\n    </Transceivers>\n    <Transducers MergeOperation=\"AddNodeTree\">\n        <Transducer TransducerName=\"ES70-7C\" TransducerSerialNumber=\"116\" TransducerCustomName=\"ES70-7C Serial No: 116\" TransducerMounting=\"HullMounted\" TransducerOffsetX=\"0\" TransducerOffsetY=\"0\" TransducerOffsetZ=\"0\" TransducerAlphaX=\"0\" TransducerAlphaY=\"0\" TransducerAlphaZ=\"0\" />\n        <Transducer TransducerName=\"ES120-7C\" TransducerSerialNumber=\"1808\" TransducerCustomName=\"ES120-7C Serial No: 1808\" TransducerMounting=\"HullMounted\" TransducerOffsetX=\"0\" TransducerOffsetY=\"0\" TransducerOffsetZ=\"0\" TransducerAlphaX=\"0\" TransducerAlphaY=\"0\" TransducerAlphaZ=\"0\" />\n        <Transducer TransducerName=\"ES200-7C\" TransducerSerialNumber=\"213\" TransducerCustomName=\"ES200-7C Serial No: 213\" TransducerMounting=\"HullMounted\" TransducerOffsetX=\"0\" TransducerOffsetY=\"0\" TransducerOffsetZ=\"0\" TransducerAlphaX=\"0\" TransducerAlphaY=\"0\" TransducerAlphaZ=\"0\" />\n    </Transducers>\n    <ConfiguredSensors MergeOperation=\"AddNodeTree\">\n        <Sensor Name=\"GPS From Serial Port 5\" Type=\"GPS\" Port=\"Serial Port 5\" TalkerID=\"\" X=\"0\" Y=\"0\" Z=\"0\" AngleX=\"0\" AngleY=\"0\" AngleZ=\"0\" Unique=\"0\" Timeout=\"20\">\n            <Telegram Name=\"GLL from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"GLL\" SubscriptionPath=\"GPS From Serial Port 5@GPS.Geographical.Position\" Enabled=\"1\">\n                <Value Name=\"Latitude\" Priority=\"1\" />\n                <Value Name=\"Longitude\" Priority=\"1\" />\n            </Telegram>\n            <Telegram Name=\"GGA from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"GGA\" SubscriptionPath=\"GPS From Serial Port 5@GPS.Global.Position\" Enabled=\"1\">\n                <Value Name=\"Latitude\" Priority=\"2\" />\n                <Value Name=\"Longitude\" Priority=\"2\" />\n            </Telegram>\n            <Telegram Name=\"GGK from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"GGK\" SubscriptionPath=\"GPS From Serial Port 5@GPS.GGK.Position\" Enabled=\"1\">\n                <Value Name=\"Latitude\" Priority=\"3\" />\n                <Value Name=\"Longitude\" Priority=\"3\" />\n            </Telegram>\n            <Telegram Name=\"PTNLGGK from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"PTNLGGK\" SubscriptionPath=\"GPS From Serial Port 5@GPS.PTNLGGK.Position\" Enabled=\"1\">\n                <Value Name=\"Latitude\" Priority=\"4\" />\n                <Value Name=\"Longitude\" Priority=\"4\" />\n            </Telegram>\n            <Telegram Name=\"RMC from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"RMC\" SubscriptionPath=\"GPS From Serial Port 5@GPS.Specific.PositionSpeedCourse\" Enabled=\"1\">\n                <Value Name=\"Latitude\" Priority=\"5\" />\n                <Value Name=\"Longitude\" Priority=\"5\" />\n                <Value Name=\"Course\" Priority=\"1\" />\n                <Value Name=\"Speed\" Priority=\"1\" />\n            </Telegram>\n            <Telegram Name=\"VTG from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"VTG\" SubscriptionPath=\"GPS From Serial Port 5@GPS.Ground\" Enabled=\"1\">\n                <Value Name=\"Course\" Priority=\"2\" />\n                <Value Name=\"CourseNotUsedMagnetic\" Priority=\"1\" />\n                <Value Name=\"Speed\" Priority=\"2\" />\n            </Telegram>\n            <Telegram Name=\"ZDA from GPS From Serial Port 5\" SensorType=\"GPS\" Type=\"ZDA\" SubscriptionPath=\"GPS From Serial Port 5@GPS.TimeInfo\" Enabled=\"1\">\n                <Value Name=\"TimeInfo\" Priority=\"1\" />\n            </Telegram>\n        </Sensor>\n    </ConfiguredSensors>\n</Configuration>" ;
  data:

   frequency_nominal = 120000, 200000, 70000 ;

   sa_correction =
  0, 0, 0, 0, -0.08,
  0, 0, 0, 0, -0.02,
  0, 0, 0, -0.02, 0 ;

   gain_correction =
  27, 27, 27, 27, 27.12,
  26, 26, 26, 26, 26.84,
  27, 27, 27, 28.88, 27 ;

   pulse_length =
  6.4e-05, 0.000128, 0.000256, 0.000512, 0.001024,
  6.4e-05, 0.000128, 0.000256, 0.000512, 0.001024,
  0.000128, 0.000256, 0.000512, 0.001024, 0.002048 ;

   channel = "WBT 150013-15 ES120-7C_ES", "WBT 545612-15 ES200-7C_ES", 
      "WBT 549762-15 ES70-7C_ES" ;

   pulse_length_bin = 0, 1, 2, 3, 4 ;

   impedance_transceiver = 5400, 5400, 5400 ;

   fs_receiver = 1500000, 1500000, 1500000 ;

   transceiver_type = "WBT", "WBT", "WBT" ;
  } // group Vendor_specific
}
